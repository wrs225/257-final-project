

module comparator_latch #
(
  parameter n_to_response_time = -1038,
  parameter p_to_response_time = -1020,
  parameter const_response_time = 1285,
  parameter n_to_tau = -1248,
  parameter p_to_tau = 1037,
  parameter const_tau = 1042,
  parameter n_to_response_time_lh = -1752,
  parameter p_to_response_time_lh = -1006,
  parameter const_response_time_lh = 1185,
  parameter n_to_tau_lh = 1131,
  parameter p_to_tau_lh = -1115,
  parameter const_tau_lh = 1529
)
(
  input clk,
  input reset,
  input sys_clk,
  input [10-1:0] n,
  input [10-1:0] p,
  output [10-1:0] out
);

  reg [17-1:0] state_cycle_counter;
  reg [1-1:0] prev_sys_clk;
  reg [35-1:0] o;
  wire [32-1:0] wait_time;
  wire [51-1:0] tau;
  wire [36-1:0] dvdt;
  wire [32-1:0] wait_time_lh;
  wire [59-1:0] tau_lh;
  wire [37-1:0] dodt;
  reg [32-1:0] fsm;
  localparam fsm_init = 0;
  wire [35-1:0] padr_0;
  wire [20-1:0] padr_bits_1;
  assign padr_bits_1 = 0;
  wire [21-1:0] truncR_2;
  wire [21-1:0] padl_3;
  wire [19-1:0] padl_bits_4;
  wire [1-1:0] toSInt_5;
  assign toSInt_5 = 0;
  wire [19-1:0] toSInt_imm_6;
  wire [18-1:0] const_7;
  assign const_7 = 18'd216268;
  assign toSInt_imm_6 = { toSInt_5, const_7 };
  assign padl_bits_4 = toSInt_imm_6;
  assign padl_3 = { { 2{ padl_bits_4[18] } }, padl_bits_4 };
  assign truncR_2 = padl_3;
  wire [15-1:0] truncR_shift_8;
  assign truncR_shift_8 = truncR_2 >>> 6;
  wire [15-1:0] truncR_imm_9;
  assign truncR_imm_9 = (truncR_2[20])? truncR_shift_8[14:0] : truncR_2[20:6];
  assign padr_0 = { truncR_imm_9, padr_bits_1 };
  wire [13-1:0] truncR_10;
  wire [14-1:0] truncval_11;
  wire [15-1:0] toUsInt_12;
  wire [35-1:0] truncR_13;
  assign truncR_13 = o;
  wire [15-1:0] truncR_shift_14;
  assign truncR_shift_14 = truncR_13 >>> 20;
  wire [15-1:0] truncR_imm_15;
  assign truncR_imm_15 = (truncR_13[34])? truncR_shift_14[14:0] : truncR_13[34:20];
  assign toUsInt_12 = truncR_imm_15;
  assign truncval_11 = toUsInt_12[11:0];
  assign truncR_10 = truncval_11[12:0];
  wire [32-1:0] padl_16;
  wire [18-1:0] padl_bits_17;
  wire [28-1:0] truncR_18;
  wire [28-1:0] padl_19;
  wire [13-1:0] padl_bits_20;
  wire [79-1:0] truncR_21;
  wire [146-1:0] truncval_22;
  wire [146-1:0] padl_23;
  wire [81-1:0] padl_bits_24;
  wire [81-1:0] padl_25;
  wire [48-1:0] padl_bits_26;
  wire [98-1:0] truncR_27;
  wire [105-1:0] truncval_28;
  wire [105-1:0] padl_29;
  wire [52-1:0] padl_bits_30;
  wire [52-1:0] padr_31;
  wire [41-1:0] padr_bits_32;
  assign padr_bits_32 = 0;
  wire [1-1:0] toSInt_33;
  assign toSInt_33 = 0;
  wire [11-1:0] toSInt_imm_34;
  assign toSInt_imm_34 = { toSInt_33, n };
  assign padr_31 = { toSInt_imm_34, padr_bits_32 };
  assign padl_bits_30 = padr_31;
  assign padl_29 = { { 53{ padl_bits_30[51] } }, padl_bits_30 };
  wire [105-1:0] padl_35;
  wire [52-1:0] padl_bits_36;
  wire [52-1:0] padl_37;
  wire [50-1:0] padl_bits_38;
  wire [50-1:0] param_39;
  assign param_39 = n_to_response_time;
  assign padl_bits_38 = param_39;
  assign padl_37 = { { 2{ padl_bits_38[49] } }, padl_bits_38 };
  assign padl_bits_36 = padl_37;
  assign padl_35 = { { 53{ padl_bits_36[51] } }, padl_bits_36 };
  assign truncval_28 = padl_29 * padl_35;
  wire [98-1:0] truncval_imm_40;
  assign truncval_imm_40 = { truncval_28[104], truncval_28[96:0] };
  assign truncR_27 = truncval_imm_40;
  wire [48-1:0] truncR_shift_41;
  assign truncR_shift_41 = truncR_27 >>> 50;
  wire [48-1:0] truncR_imm_42;
  assign truncR_imm_42 = (truncR_27[97])? truncR_shift_41[47:0] : truncR_27[97:50];
  wire [48-1:0] padr_43;
  wire [2-1:0] padr_bits_44;
  assign padr_bits_44 = 0;
  wire [94-1:0] truncR_45;
  wire [101-1:0] truncval_46;
  wire [101-1:0] padl_47;
  wire [50-1:0] padl_bits_48;
  wire [50-1:0] padr_49;
  wire [39-1:0] padr_bits_50;
  assign padr_bits_50 = 0;
  wire [1-1:0] toSInt_51;
  assign toSInt_51 = 0;
  wire [11-1:0] toSInt_imm_52;
  assign toSInt_imm_52 = { toSInt_51, p };
  assign padr_49 = { toSInt_imm_52, padr_bits_50 };
  assign padl_bits_48 = padr_49;
  assign padl_47 = { { 51{ padl_bits_48[49] } }, padl_bits_48 };
  wire [101-1:0] padl_53;
  wire [50-1:0] padl_bits_54;
  wire [50-1:0] padl_55;
  wire [48-1:0] padl_bits_56;
  wire [48-1:0] param_57;
  assign param_57 = p_to_response_time;
  assign padl_bits_56 = param_57;
  assign padl_55 = { { 2{ padl_bits_56[47] } }, padl_bits_56 };
  assign padl_bits_54 = padl_55;
  assign padl_53 = { { 51{ padl_bits_54[49] } }, padl_bits_54 };
  assign truncval_46 = padl_47 * padl_53;
  wire [94-1:0] truncval_imm_58;
  assign truncval_imm_58 = { truncval_46[100], truncval_46[92:0] };
  assign truncR_45 = truncval_imm_58;
  wire [46-1:0] truncR_shift_59;
  assign truncR_shift_59 = truncR_45 >>> 48;
  wire [46-1:0] truncR_imm_60;
  assign truncR_imm_60 = (truncR_45[93])? truncR_shift_59[45:0] : truncR_45[93:48];
  assign padr_43 = { truncR_imm_60, padr_bits_44 };
  wire [48-1:0] padr_61;
  wire [4-1:0] padr_bits_62;
  assign padr_bits_62 = 0;
  wire [44-1:0] padl_63;
  wire [43-1:0] padl_bits_64;
  wire [1-1:0] toSInt_65;
  assign toSInt_65 = 0;
  wire [43-1:0] toSInt_imm_66;
  wire [42-1:0] param_67;
  assign param_67 = const_response_time;
  assign toSInt_imm_66 = { toSInt_65, param_67 };
  assign padl_bits_64 = toSInt_imm_66;
  assign padl_63 = { { 1{ padl_bits_64[42] } }, padl_bits_64 };
  assign padr_61 = { padl_63, padr_bits_62 };
  assign padl_bits_26 = truncR_imm_42 + padr_43 + padr_61;
  assign padl_25 = { { 33{ padl_bits_26[47] } }, padl_bits_26 };
  assign padl_bits_24 = padl_25;
  assign padl_23 = { { 65{ padl_bits_24[80] } }, padl_bits_24 };
  wire [146-1:0] padl_68;
  wire [81-1:0] padl_bits_69;
  wire [81-1:0] padr_70;
  wire [46-1:0] padr_bits_71;
  assign padr_bits_71 = 0;
  wire [1-1:0] toSInt_72;
  assign toSInt_72 = 0;
  wire [35-1:0] toSInt_imm_73;
  wire [34-1:0] const_74;
  assign const_74 = 34'd152587;
  assign toSInt_imm_73 = { toSInt_72, const_74 };
  assign padr_70 = { toSInt_imm_73, padr_bits_71 };
  assign padl_bits_69 = padr_70;
  assign padl_68 = { { 65{ padl_bits_69[80] } }, padl_bits_69 };
  assign truncval_22 = padl_23 * padl_68;
  assign truncR_21 = truncval_22[78:0];
  assign padl_bits_20 = truncR_21[78:66];
  wire [15-1:0] padl_bits_zero_75;
  assign padl_bits_zero_75 = 0;
  assign padl_19 = { padl_bits_zero_75, padl_bits_20 };
  assign truncR_18 = padl_19;
  assign padl_bits_17 = truncR_18[27:10];
  wire [14-1:0] padl_bits_zero_76;
  assign padl_bits_zero_76 = 0;
  assign padl_16 = { padl_bits_zero_76, padl_bits_17 };
  assign wait_time = padl_16;
  wire [35-1:0] padr_77;
  wire [20-1:0] padr_bits_78;
  assign padr_bits_78 = 0;
  wire [21-1:0] truncR_79;
  wire [21-1:0] padl_80;
  wire [19-1:0] padl_bits_81;
  wire [1-1:0] toSInt_82;
  assign toSInt_82 = 0;
  wire [19-1:0] toSInt_imm_83;
  wire [18-1:0] const_84;
  assign const_84 = 18'd216268;
  assign toSInt_imm_83 = { toSInt_82, const_84 };
  assign padl_bits_81 = toSInt_imm_83;
  assign padl_80 = { { 2{ padl_bits_81[18] } }, padl_bits_81 };
  assign truncR_79 = padl_80;
  wire [15-1:0] truncR_shift_85;
  assign truncR_shift_85 = truncR_79 >>> 6;
  wire [15-1:0] truncR_imm_86;
  assign truncR_imm_86 = (truncR_79[20])? truncR_shift_85[14:0] : truncR_79[20:6];
  assign padr_77 = { truncR_imm_86, padr_bits_78 };
  wire [13-1:0] truncR_87;
  wire [14-1:0] truncval_88;
  wire [15-1:0] toUsInt_89;
  wire [35-1:0] truncR_90;
  assign truncR_90 = o;
  wire [15-1:0] truncR_shift_91;
  assign truncR_shift_91 = truncR_90 >>> 20;
  wire [15-1:0] truncR_imm_92;
  assign truncR_imm_92 = (truncR_90[34])? truncR_shift_91[14:0] : truncR_90[34:20];
  assign toUsInt_89 = truncR_imm_92;
  assign truncval_88 = toUsInt_89[11:0];
  assign truncR_87 = truncval_88[12:0];
  wire [51-1:0] padr_93;
  wire [10-1:0] padr_bits_94;
  assign padr_bits_94 = 0;
  wire [42-1:0] truncval_95;
  wire [43-1:0] toUsInt_96;
  wire [43-1:0] padr_97;
  wire [1-1:0] padr_bits_98;
  assign padr_bits_98 = 0;
  wire [88-1:0] truncR_99;
  wire [95-1:0] truncval_100;
  wire [95-1:0] padl_101;
  wire [47-1:0] padl_bits_102;
  wire [47-1:0] padr_103;
  wire [36-1:0] padr_bits_104;
  assign padr_bits_104 = 0;
  wire [1-1:0] toSInt_105;
  assign toSInt_105 = 0;
  wire [11-1:0] toSInt_imm_106;
  assign toSInt_imm_106 = { toSInt_105, n };
  assign padr_103 = { toSInt_imm_106, padr_bits_104 };
  assign padl_bits_102 = padr_103;
  assign padl_101 = { { 48{ padl_bits_102[46] } }, padl_bits_102 };
  wire [95-1:0] padl_107;
  wire [47-1:0] padl_bits_108;
  wire [47-1:0] padl_109;
  wire [45-1:0] padl_bits_110;
  wire [45-1:0] param_111;
  assign param_111 = n_to_tau;
  assign padl_bits_110 = param_111;
  assign padl_109 = { { 2{ padl_bits_110[44] } }, padl_bits_110 };
  assign padl_bits_108 = padl_109;
  assign padl_107 = { { 48{ padl_bits_108[46] } }, padl_bits_108 };
  assign truncval_100 = padl_101 * padl_107;
  wire [88-1:0] truncval_imm_112;
  assign truncval_imm_112 = { truncval_100[94], truncval_100[86:0] };
  assign truncR_99 = truncval_imm_112;
  wire [42-1:0] truncR_shift_113;
  assign truncR_shift_113 = truncR_99 >>> 46;
  wire [42-1:0] truncR_imm_114;
  assign truncR_imm_114 = (truncR_99[87])? truncR_shift_113[41:0] : truncR_99[87:46];
  assign padr_97 = { truncR_imm_114, padr_bits_98 };
  wire [43-1:0] padl_115;
  wire [42-1:0] padl_bits_116;
  wire [1-1:0] toSInt_117;
  assign toSInt_117 = 0;
  wire [42-1:0] toSInt_imm_118;
  wire [86-1:0] truncR_119;
  wire [92-1:0] truncval_120;
  wire [92-1:0] padl_121;
  wire [46-1:0] padl_bits_122;
  wire [46-1:0] padr_123;
  wire [36-1:0] padr_bits_124;
  assign padr_bits_124 = 0;
  assign padr_123 = { p, padr_bits_124 };
  assign padl_bits_122 = padr_123;
  wire [46-1:0] padl_bits_zero_125;
  assign padl_bits_zero_125 = 0;
  assign padl_121 = { padl_bits_zero_125, padl_bits_122 };
  wire [92-1:0] padl_126;
  wire [46-1:0] padl_bits_127;
  wire [46-1:0] padl_128;
  wire [43-1:0] padl_bits_129;
  wire [43-1:0] param_130;
  assign param_130 = p_to_tau;
  assign padl_bits_129 = param_130;
  wire [3-1:0] padl_bits_zero_131;
  assign padl_bits_zero_131 = 0;
  assign padl_128 = { padl_bits_zero_131, padl_bits_129 };
  assign padl_bits_127 = padl_128;
  wire [46-1:0] padl_bits_zero_132;
  assign padl_bits_zero_132 = 0;
  assign padl_126 = { padl_bits_zero_132, padl_bits_127 };
  assign truncval_120 = padl_121 * padl_126;
  assign truncR_119 = truncval_120[85:0];
  assign toSInt_imm_118 = { toSInt_117, truncR_119[85:45] };
  assign padl_bits_116 = toSInt_imm_118;
  assign padl_115 = { { 1{ padl_bits_116[41] } }, padl_bits_116 };
  wire [43-1:0] padl_133;
  wire [42-1:0] padl_bits_134;
  wire [1-1:0] toSInt_135;
  assign toSInt_135 = 0;
  wire [42-1:0] toSInt_imm_136;
  wire [41-1:0] param_137;
  assign param_137 = const_tau;
  assign toSInt_imm_136 = { toSInt_135, param_137 };
  assign padl_bits_134 = toSInt_imm_136;
  assign padl_133 = { { 1{ padl_bits_134[41] } }, padl_bits_134 };
  assign toUsInt_96 = padr_97 + padl_115 + padl_133;
  assign truncval_95 = toUsInt_96[39:0];
  assign padr_93 = { truncval_95[40:0], padr_bits_94 };
  assign tau = padr_93;
  wire [13-1:0] truncR_138;
  wire [14-1:0] truncval_139;
  wire [15-1:0] toUsInt_140;
  wire [35-1:0] truncR_141;
  assign truncR_141 = o;
  wire [15-1:0] truncR_shift_142;
  assign truncR_shift_142 = truncR_141 >>> 20;
  wire [15-1:0] truncR_imm_143;
  assign truncR_imm_143 = (truncR_141[34])? truncR_shift_142[14:0] : truncR_141[34:20];
  assign toUsInt_140 = truncR_imm_143;
  assign truncval_139 = toUsInt_140[11:0];
  assign truncR_138 = truncval_139[12:0];
  wire [36-1:0] padl_144;
  wire [13-1:0] padl_bits_145;
  wire [36-1:0] truncR_146;
  wire [50-1:0] truncR_147;
  wire [83-1:0] truncval_148;
  wire [83-1:0] padl_149;
  wire [41-1:0] padl_bits_150;
  wire [41-1:0] padl_151;
  wire [12-1:0] padl_bits_152;
  wire [12-1:0] neg_imm_153;
  wire [15-1:0] truncR_154;
  wire [35-1:0] truncR_155;
  assign truncR_155 = o;
  wire [15-1:0] truncR_shift_156;
  assign truncR_shift_156 = truncR_155 >>> 20;
  wire [15-1:0] truncR_imm_157;
  assign truncR_imm_157 = (truncR_155[34])? truncR_shift_156[14:0] : truncR_155[34:20];
  assign truncR_154 = truncR_imm_157;
  wire [12-1:0] truncR_shift_158;
  assign truncR_shift_158 = truncR_154 >>> 3;
  wire [12-1:0] truncR_imm_159;
  assign truncR_imm_159 = (truncR_154[14])? truncR_shift_158[11:0] : truncR_154[14:3];
  assign neg_imm_153 = -truncR_imm_159;
  assign padl_bits_152 = neg_imm_153;
  assign padl_151 = { { 29{ padl_bits_152[11] } }, padl_bits_152 };
  assign padl_bits_150 = padl_151;
  assign padl_149 = { { 42{ padl_bits_150[40] } }, padl_bits_150 };
  wire [83-1:0] padl_160;
  wire [41-1:0] padl_bits_161;
  wire [41-1:0] padr_162;
  wire [7-1:0] padr_bits_163;
  assign padr_bits_163 = 0;
  wire [1-1:0] toSInt_164;
  assign toSInt_164 = 0;
  wire [34-1:0] toSInt_imm_165;
  wire [51-1:0] truncval_166;
  assign truncval_166 = 52'd2251799813685248 / tau;
  assign toSInt_imm_165 = { toSInt_164, truncval_166[32:0] };
  assign padr_162 = { toSInt_imm_165, padr_bits_163 };
  assign padl_bits_161 = padr_162;
  assign padl_160 = { { 42{ padl_bits_161[40] } }, padl_bits_161 };
  assign truncval_148 = padl_149 * padl_160;
  wire [50-1:0] truncval_imm_167;
  assign truncval_imm_167 = { truncval_148[82], truncval_148[48:0] };
  assign truncR_147 = truncval_imm_167;
  wire [36-1:0] truncR_shift_168;
  assign truncR_shift_168 = truncR_147 >>> 14;
  wire [36-1:0] truncR_imm_169;
  assign truncR_imm_169 = (truncR_147[49])? truncR_shift_168[35:0] : truncR_147[49:14];
  assign truncR_146 = truncR_imm_169;
  wire [13-1:0] truncR_shift_170;
  assign truncR_shift_170 = truncR_146 >>> 23;
  wire [13-1:0] truncR_imm_171;
  assign truncR_imm_171 = (truncR_146[35])? truncR_shift_170[12:0] : truncR_146[35:23];
  assign padl_bits_145 = truncR_imm_171;
  assign padl_144 = { { 23{ padl_bits_145[12] } }, padl_bits_145 };
  assign dvdt = padl_144;
  wire [35-1:0] padr_172;
  wire [20-1:0] padr_bits_173;
  assign padr_bits_173 = 0;
  wire [15-1:0] padr_174;
  wire [1-1:0] padr_bits_175;
  assign padr_bits_175 = 0;
  wire [14-1:0] padl_176;
  wire [12-1:0] padl_bits_177;
  wire [82-1:0] truncR_178;
  wire [152-1:0] truncval_179;
  wire [152-1:0] padl_180;
  wire [87-1:0] padl_bits_181;
  wire [87-1:0] padl_182;
  wire [52-1:0] padl_bits_183;
  wire [1-1:0] toSInt_184;
  assign toSInt_184 = 0;
  wire [52-1:0] toSInt_imm_185;
  wire [51-1:0] const_186;
  assign const_186 = 51'd225179;
  assign toSInt_imm_185 = { toSInt_184, const_186 };
  assign padl_bits_183 = toSInt_imm_185;
  assign padl_182 = { { 35{ padl_bits_183[51] } }, padl_bits_183 };
  assign padl_bits_181 = padl_182;
  assign padl_180 = { { 65{ padl_bits_181[86] } }, padl_bits_181 };
  wire [152-1:0] padl_187;
  wire [87-1:0] padl_bits_188;
  wire [87-1:0] padr_189;
  wire [51-1:0] padr_bits_190;
  assign padr_bits_190 = 0;
  assign padr_189 = { dvdt, padr_bits_190 };
  assign padl_bits_188 = padr_189;
  assign padl_187 = { { 65{ padl_bits_188[86] } }, padl_bits_188 };
  assign truncval_179 = padl_180 * padl_187;
  wire [82-1:0] truncval_imm_191;
  assign truncval_imm_191 = { truncval_179[151], truncval_179[80:0] };
  assign truncR_178 = truncval_imm_191;
  wire [12-1:0] truncR_shift_192;
  assign truncR_shift_192 = truncR_178 >>> 70;
  wire [12-1:0] truncR_imm_193;
  assign truncR_imm_193 = (truncR_178[81])? truncR_shift_192[11:0] : truncR_178[81:70];
  assign padl_bits_177 = truncR_imm_193;
  assign padl_176 = { { 2{ padl_bits_177[11] } }, padl_bits_177 };
  assign padr_174 = { padl_176, padr_bits_175 };
  assign padr_172 = { padr_174, padr_bits_173 };
  wire [32-1:0] padl_194;
  wire [2-1:0] padl_bits_195;
  wire [13-1:0] truncR_196;
  wire [13-1:0] padr_197;
  wire [1-1:0] padr_bits_198;
  assign padr_bits_198 = 0;
  wire [76-1:0] truncR_199;
  wire [144-1:0] truncval_200;
  wire [144-1:0] padl_201;
  wire [80-1:0] padl_bits_202;
  wire [80-1:0] padl_203;
  wire [47-1:0] padl_bits_204;
  wire [98-1:0] truncR_205;
  wire [105-1:0] truncval_206;
  wire [105-1:0] padl_207;
  wire [52-1:0] padl_bits_208;
  wire [52-1:0] padr_209;
  wire [41-1:0] padr_bits_210;
  assign padr_bits_210 = 0;
  wire [1-1:0] toSInt_211;
  assign toSInt_211 = 0;
  wire [11-1:0] toSInt_imm_212;
  assign toSInt_imm_212 = { toSInt_211, n };
  assign padr_209 = { toSInt_imm_212, padr_bits_210 };
  assign padl_bits_208 = padr_209;
  assign padl_207 = { { 53{ padl_bits_208[51] } }, padl_bits_208 };
  wire [105-1:0] padl_213;
  wire [52-1:0] padl_bits_214;
  wire [52-1:0] padl_215;
  wire [50-1:0] padl_bits_216;
  wire [50-1:0] param_217;
  assign param_217 = n_to_response_time_lh;
  assign padl_bits_216 = param_217;
  assign padl_215 = { { 2{ padl_bits_216[49] } }, padl_bits_216 };
  assign padl_bits_214 = padl_215;
  assign padl_213 = { { 53{ padl_bits_214[51] } }, padl_bits_214 };
  assign truncval_206 = padl_207 * padl_213;
  wire [98-1:0] truncval_imm_218;
  assign truncval_imm_218 = { truncval_206[104], truncval_206[96:0] };
  assign truncR_205 = truncval_imm_218;
  wire [47-1:0] truncR_shift_219;
  assign truncR_shift_219 = truncR_205 >>> 51;
  wire [47-1:0] truncR_imm_220;
  assign truncR_imm_220 = (truncR_205[97])? truncR_shift_219[46:0] : truncR_205[97:51];
  wire [47-1:0] padr_221;
  wire [1-1:0] padr_bits_222;
  assign padr_bits_222 = 0;
  wire [94-1:0] truncR_223;
  wire [101-1:0] truncval_224;
  wire [101-1:0] padl_225;
  wire [50-1:0] padl_bits_226;
  wire [50-1:0] padr_227;
  wire [39-1:0] padr_bits_228;
  assign padr_bits_228 = 0;
  wire [1-1:0] toSInt_229;
  assign toSInt_229 = 0;
  wire [11-1:0] toSInt_imm_230;
  assign toSInt_imm_230 = { toSInt_229, p };
  assign padr_227 = { toSInt_imm_230, padr_bits_228 };
  assign padl_bits_226 = padr_227;
  assign padl_225 = { { 51{ padl_bits_226[49] } }, padl_bits_226 };
  wire [101-1:0] padl_231;
  wire [50-1:0] padl_bits_232;
  wire [50-1:0] padl_233;
  wire [48-1:0] padl_bits_234;
  wire [48-1:0] param_235;
  assign param_235 = p_to_response_time_lh;
  assign padl_bits_234 = param_235;
  assign padl_233 = { { 2{ padl_bits_234[47] } }, padl_bits_234 };
  assign padl_bits_232 = padl_233;
  assign padl_231 = { { 51{ padl_bits_232[49] } }, padl_bits_232 };
  assign truncval_224 = padl_225 * padl_231;
  wire [94-1:0] truncval_imm_236;
  assign truncval_imm_236 = { truncval_224[100], truncval_224[92:0] };
  assign truncR_223 = truncval_imm_236;
  wire [46-1:0] truncR_shift_237;
  assign truncR_shift_237 = truncR_223 >>> 48;
  wire [46-1:0] truncR_imm_238;
  assign truncR_imm_238 = (truncR_223[93])? truncR_shift_237[45:0] : truncR_223[93:48];
  assign padr_221 = { truncR_imm_238, padr_bits_222 };
  wire [47-1:0] padr_239;
  wire [2-1:0] padr_bits_240;
  assign padr_bits_240 = 0;
  wire [45-1:0] padl_241;
  wire [44-1:0] padl_bits_242;
  wire [1-1:0] toSInt_243;
  assign toSInt_243 = 0;
  wire [44-1:0] toSInt_imm_244;
  wire [43-1:0] param_245;
  assign param_245 = const_response_time_lh;
  assign toSInt_imm_244 = { toSInt_243, param_245 };
  assign padl_bits_242 = toSInt_imm_244;
  assign padl_241 = { { 1{ padl_bits_242[43] } }, padl_bits_242 };
  assign padr_239 = { padl_241, padr_bits_240 };
  assign padl_bits_204 = truncR_imm_220 + padr_221 + padr_239;
  assign padl_203 = { { 33{ padl_bits_204[46] } }, padl_bits_204 };
  assign padl_bits_202 = padl_203;
  assign padl_201 = { { 64{ padl_bits_202[79] } }, padl_bits_202 };
  wire [144-1:0] padl_246;
  wire [80-1:0] padl_bits_247;
  wire [80-1:0] padr_248;
  wire [45-1:0] padr_bits_249;
  assign padr_bits_249 = 0;
  wire [1-1:0] toSInt_250;
  assign toSInt_250 = 0;
  wire [35-1:0] toSInt_imm_251;
  wire [34-1:0] const_252;
  assign const_252 = 34'd152587;
  assign toSInt_imm_251 = { toSInt_250, const_252 };
  assign padr_248 = { toSInt_imm_251, padr_bits_249 };
  assign padl_bits_247 = padr_248;
  assign padl_246 = { { 64{ padl_bits_247[79] } }, padl_bits_247 };
  assign truncval_200 = padl_201 * padl_246;
  assign truncR_199 = truncval_200[75:0];
  assign padr_197 = { truncR_199[75:64], padr_bits_198 };
  assign truncR_196 = padr_197;
  assign padl_bits_195 = truncR_196[12:11];
  wire [30-1:0] padl_bits_zero_253;
  assign padl_bits_zero_253 = 0;
  assign padl_194 = { padl_bits_zero_253, padl_bits_195 };
  assign wait_time_lh = padl_194;
  wire [35-1:0] padr_254;
  wire [20-1:0] padr_bits_255;
  assign padr_bits_255 = 0;
  wire [32-1:0] truncR_256;
  wire [32-1:0] padl_257;
  wire [28-1:0] padl_bits_258;
  wire [1-1:0] toSInt_259;
  assign toSInt_259 = 0;
  wire [28-1:0] toSInt_imm_260;
  wire [27-1:0] const_261;
  assign const_261 = 27'd134217;
  assign toSInt_imm_260 = { toSInt_259, const_261 };
  assign padl_bits_258 = toSInt_imm_260;
  assign padl_257 = { { 4{ padl_bits_258[27] } }, padl_bits_258 };
  assign truncR_256 = padl_257;
  wire [15-1:0] truncR_shift_262;
  assign truncR_shift_262 = truncR_256 >>> 17;
  wire [15-1:0] truncR_imm_263;
  assign truncR_imm_263 = (truncR_256[31])? truncR_shift_262[14:0] : truncR_256[31:17];
  assign padr_254 = { truncR_imm_263, padr_bits_255 };
  wire [13-1:0] truncR_264;
  wire [14-1:0] truncval_265;
  wire [15-1:0] toUsInt_266;
  wire [35-1:0] truncR_267;
  assign truncR_267 = o;
  wire [15-1:0] truncR_shift_268;
  assign truncR_shift_268 = truncR_267 >>> 20;
  wire [15-1:0] truncR_imm_269;
  assign truncR_imm_269 = (truncR_267[34])? truncR_shift_268[14:0] : truncR_267[34:20];
  assign toUsInt_266 = truncR_imm_269;
  assign truncval_265 = toUsInt_266[11:0];
  assign truncR_264 = truncval_265[12:0];
  wire [59-1:0] padr_270;
  wire [14-1:0] padr_bits_271;
  assign padr_bits_271 = 0;
  wire [46-1:0] truncval_272;
  wire [47-1:0] toUsInt_273;
  wire [47-1:0] padr_274;
  wire [3-1:0] padr_bits_275;
  assign padr_bits_275 = 0;
  wire [44-1:0] padl_276;
  wire [43-1:0] padl_bits_277;
  wire [1-1:0] toSInt_278;
  assign toSInt_278 = 0;
  wire [43-1:0] toSInt_imm_279;
  wire [88-1:0] truncR_280;
  wire [94-1:0] truncval_281;
  wire [94-1:0] padl_282;
  wire [47-1:0] padl_bits_283;
  wire [47-1:0] padr_284;
  wire [37-1:0] padr_bits_285;
  assign padr_bits_285 = 0;
  assign padr_284 = { n, padr_bits_285 };
  assign padl_bits_283 = padr_284;
  wire [47-1:0] padl_bits_zero_286;
  assign padl_bits_zero_286 = 0;
  assign padl_282 = { padl_bits_zero_286, padl_bits_283 };
  wire [94-1:0] padl_287;
  wire [47-1:0] padl_bits_288;
  wire [47-1:0] padl_289;
  wire [44-1:0] padl_bits_290;
  wire [44-1:0] param_291;
  assign param_291 = n_to_tau_lh;
  assign padl_bits_290 = param_291;
  wire [3-1:0] padl_bits_zero_292;
  assign padl_bits_zero_292 = 0;
  assign padl_289 = { padl_bits_zero_292, padl_bits_290 };
  assign padl_bits_288 = padl_289;
  wire [47-1:0] padl_bits_zero_293;
  assign padl_bits_zero_293 = 0;
  assign padl_287 = { padl_bits_zero_293, padl_bits_288 };
  assign truncval_281 = padl_282 * padl_287;
  assign truncR_280 = truncval_281[87:0];
  assign toSInt_imm_279 = { toSInt_278, truncR_280[87:46] };
  assign padl_bits_277 = toSInt_imm_279;
  assign padl_276 = { { 1{ padl_bits_277[42] } }, padl_bits_277 };
  assign padr_274 = { padl_276, padr_bits_275 };
  wire [96-1:0] truncR_294;
  wire [103-1:0] truncval_295;
  wire [103-1:0] padl_296;
  wire [51-1:0] padl_bits_297;
  wire [51-1:0] padr_298;
  wire [40-1:0] padr_bits_299;
  assign padr_bits_299 = 0;
  wire [1-1:0] toSInt_300;
  assign toSInt_300 = 0;
  wire [11-1:0] toSInt_imm_301;
  assign toSInt_imm_301 = { toSInt_300, p };
  assign padr_298 = { toSInt_imm_301, padr_bits_299 };
  assign padl_bits_297 = padr_298;
  assign padl_296 = { { 52{ padl_bits_297[50] } }, padl_bits_297 };
  wire [103-1:0] padl_302;
  wire [51-1:0] padl_bits_303;
  wire [51-1:0] padl_304;
  wire [49-1:0] padl_bits_305;
  wire [49-1:0] param_306;
  assign param_306 = p_to_tau_lh;
  assign padl_bits_305 = param_306;
  assign padl_304 = { { 2{ padl_bits_305[48] } }, padl_bits_305 };
  assign padl_bits_303 = padl_304;
  assign padl_302 = { { 52{ padl_bits_303[50] } }, padl_bits_303 };
  assign truncval_295 = padl_296 * padl_302;
  wire [96-1:0] truncval_imm_307;
  assign truncval_imm_307 = { truncval_295[102], truncval_295[94:0] };
  assign truncR_294 = truncval_imm_307;
  wire [47-1:0] truncR_shift_308;
  assign truncR_shift_308 = truncR_294 >>> 49;
  wire [47-1:0] truncR_imm_309;
  assign truncR_imm_309 = (truncR_294[95])? truncR_shift_308[46:0] : truncR_294[95:49];
  wire [47-1:0] padr_310;
  wire [2-1:0] padr_bits_311;
  assign padr_bits_311 = 0;
  wire [45-1:0] padl_312;
  wire [44-1:0] padl_bits_313;
  wire [1-1:0] toSInt_314;
  assign toSInt_314 = 0;
  wire [44-1:0] toSInt_imm_315;
  wire [43-1:0] param_316;
  assign param_316 = const_tau_lh;
  assign toSInt_imm_315 = { toSInt_314, param_316 };
  assign padl_bits_313 = toSInt_imm_315;
  assign padl_312 = { { 1{ padl_bits_313[43] } }, padl_bits_313 };
  assign padr_310 = { padl_312, padr_bits_311 };
  assign toUsInt_273 = padr_274 + truncR_imm_309 + padr_310;
  assign truncval_272 = toUsInt_273[43:0];
  assign padr_270 = { truncval_272[44:0], padr_bits_271 };
  assign tau_lh = padr_270;
  wire [33-1:0] truncR_317;
  wire [34-1:0] truncval_318;
  wire [35-1:0] toUsInt_319;
  assign toUsInt_319 = o;
  assign truncval_318 = toUsInt_319[31:0];
  assign truncR_317 = truncval_318[32:0];
  wire [37-1:0] padl_320;
  wire [13-1:0] padl_bits_321;
  wire [37-1:0] truncR_322;
  wire [97-1:0] truncR_323;
  wire [129-1:0] truncval_324;
  wire [129-1:0] padl_325;
  wire [64-1:0] padl_bits_326;
  wire [64-1:0] padl_327;
  wire [35-1:0] padl_bits_328;
  wire [35-1:0] padr_329;
  wire [14-1:0] padr_bits_330;
  assign padr_bits_330 = 0;
  wire [21-1:0] padl_331;
  wire [19-1:0] padl_bits_332;
  wire [1-1:0] toSInt_333;
  assign toSInt_333 = 0;
  wire [19-1:0] toSInt_imm_334;
  wire [18-1:0] const_335;
  assign const_335 = 18'd216268;
  assign toSInt_imm_334 = { toSInt_333, const_335 };
  assign padl_bits_332 = toSInt_imm_334;
  assign padl_331 = { { 2{ padl_bits_332[18] } }, padl_bits_332 };
  assign padr_329 = { padl_331, padr_bits_330 };
  assign padl_bits_328 = padr_329 - o;
  assign padl_327 = { { 29{ padl_bits_328[34] } }, padl_bits_328 };
  assign padl_bits_326 = padl_327;
  assign padl_325 = { { 65{ padl_bits_326[63] } }, padl_bits_326 };
  wire [129-1:0] padl_336;
  wire [64-1:0] padl_bits_337;
  wire [64-1:0] padr_338;
  wire [30-1:0] padr_bits_339;
  assign padr_bits_339 = 0;
  wire [1-1:0] toSInt_340;
  assign toSInt_340 = 0;
  wire [34-1:0] toSInt_imm_341;
  wire [59-1:0] truncval_342;
  assign truncval_342 = 60'd576460752303423488 / tau_lh;
  assign toSInt_imm_341 = { toSInt_340, truncval_342[32:0] };
  assign padr_338 = { toSInt_imm_341, padr_bits_339 };
  assign padl_bits_337 = padr_338;
  assign padl_336 = { { 65{ padl_bits_337[63] } }, padl_bits_337 };
  assign truncval_324 = padl_325 * padl_336;
  wire [97-1:0] truncval_imm_343;
  assign truncval_imm_343 = { truncval_324[128], truncval_324[95:0] };
  assign truncR_323 = truncval_imm_343;
  wire [37-1:0] truncR_shift_344;
  assign truncR_shift_344 = truncR_323 >>> 60;
  wire [37-1:0] truncR_imm_345;
  assign truncR_imm_345 = (truncR_323[96])? truncR_shift_344[36:0] : truncR_323[96:60];
  assign truncR_322 = truncR_imm_345;
  wire [13-1:0] truncR_shift_346;
  assign truncR_shift_346 = truncR_322 >>> 24;
  wire [13-1:0] truncR_imm_347;
  assign truncR_imm_347 = (truncR_322[36])? truncR_shift_346[12:0] : truncR_322[36:24];
  assign padl_bits_321 = truncR_imm_347;
  assign padl_320 = { { 24{ padl_bits_321[12] } }, padl_bits_321 };
  assign dodt = padl_320;
  wire [35-1:0] padr_348;
  wire [21-1:0] padr_bits_349;
  assign padr_bits_349 = 0;
  wire [14-1:0] padl_350;
  wire [12-1:0] padl_bits_351;
  wire [81-1:0] truncR_352;
  wire [153-1:0] truncval_353;
  wire [153-1:0] padl_354;
  wire [88-1:0] padl_bits_355;
  wire [88-1:0] padl_356;
  wire [52-1:0] padl_bits_357;
  wire [1-1:0] toSInt_358;
  assign toSInt_358 = 0;
  wire [52-1:0] toSInt_imm_359;
  wire [51-1:0] const_360;
  assign const_360 = 51'd225179;
  assign toSInt_imm_359 = { toSInt_358, const_360 };
  assign padl_bits_357 = toSInt_imm_359;
  assign padl_356 = { { 36{ padl_bits_357[51] } }, padl_bits_357 };
  assign padl_bits_355 = padl_356;
  assign padl_354 = { { 65{ padl_bits_355[87] } }, padl_bits_355 };
  wire [153-1:0] padl_361;
  wire [88-1:0] padl_bits_362;
  wire [88-1:0] padr_363;
  wire [51-1:0] padr_bits_364;
  assign padr_bits_364 = 0;
  assign padr_363 = { dodt, padr_bits_364 };
  assign padl_bits_362 = padr_363;
  assign padl_361 = { { 65{ padl_bits_362[87] } }, padl_bits_362 };
  assign truncval_353 = padl_354 * padl_361;
  wire [81-1:0] truncval_imm_365;
  assign truncval_imm_365 = { truncval_353[152], truncval_353[79:0] };
  assign truncR_352 = truncval_imm_365;
  wire [12-1:0] truncR_shift_366;
  assign truncR_shift_366 = truncR_352 >>> 69;
  wire [12-1:0] truncR_imm_367;
  assign truncR_imm_367 = (truncR_352[80])? truncR_shift_366[11:0] : truncR_352[80:69];
  assign padl_bits_351 = truncR_imm_367;
  assign padl_350 = { { 2{ padl_bits_351[11] } }, padl_bits_351 };
  assign padr_348 = { padl_350, padr_bits_349 };
  assign out = (fsm == 0)? truncR_10[12:3] : truncR_87[12:3];

  always @(posedge clk) begin
    prev_sys_clk <= sys_clk;
  end

  localparam fsm_1 = 1;
  localparam fsm_2 = 2;
  localparam fsm_3 = 3;
  localparam fsm_4 = 4;

  always @(posedge clk) begin
    if(reset) begin
      fsm <= fsm_init;
    end else begin
      case(fsm)
        fsm_init: begin
          if(reset) begin
            o <= 35'd3543348019;
          end else begin
            o <= padr_0;
          end
          if(~prev_sys_clk & sys_clk & ((n > p) & (n <= 10'd512))) begin
            fsm <= fsm_1;
          end 
        end
        fsm_1: begin
          if(reset) begin
            o <= 35'd3543348019;
          end else begin
            o <= padr_77;
          end
          if(state_cycle_counter > wait_time) begin
            state_cycle_counter <= 0;
          end else begin
            state_cycle_counter <= state_cycle_counter + 1;
          end
          if(state_cycle_counter > wait_time) begin
            fsm <= fsm_2;
          end 
        end
        fsm_2: begin
          if(reset) begin
            o <= 35'd3543348019;
          end else begin
            o <= o + padr_172;
          end
          if(prev_sys_clk & ~sys_clk) begin
            fsm <= fsm_3;
          end 
        end
        fsm_3: begin
          if(reset) begin
            o <= 35'd3543348019;
          end else begin
            o <= padr_254;
          end
          if(state_cycle_counter > wait_time_lh) begin
            state_cycle_counter <= 0;
          end else begin
            state_cycle_counter <= state_cycle_counter + 1;
          end
          if(state_cycle_counter > wait_time_lh) begin
            fsm <= fsm_4;
          end 
        end
        fsm_4: begin
          if(reset) begin
            o <= 35'd3543348019;
          end else begin
            o <= o + padr_348;
          end
          if((o > 35'd3532610600) & (o <= 35'd17179869184)) begin
            fsm <= fsm_init;
          end 
        end
      endcase
    end
  end


endmodule

