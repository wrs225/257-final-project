

module comparator_latch #
(
  parameter n_to_response_time = -1038,
  parameter p_to_response_time = -1020,
  parameter const_response_time = 1285,
  parameter n_to_tau = -1248,
  parameter p_to_tau = 1037,
  parameter const_tau = 1042,
  parameter n_to_response_time_lh = -1752,
  parameter p_to_response_time_lh = -1006,
  parameter const_response_time_lh = 1185,
  parameter n_to_tau_lh = 1131,
  parameter p_to_tau_lh = -1115,
  parameter const_tau_lh = 1529
)
(
  input clk,
  input reset,
  input sys_clk,
  input [10-1:0] n,
  input [10-1:0] p,
  output [10-1:0] out
);

  reg [17-1:0] state_cycle_counter;
  reg [1-1:0] prev_sys_clk;
  reg [35-1:0] o;
  wire [32-1:0] wait_time;
  wire [51-1:0] tau;
  wire [36-1:0] dvdt;
  wire [32-1:0] wait_time_lh;
  wire [59-1:0] tau_lh;
  wire [37-1:0] dodt;
  reg [32-1:0] fsm;
  localparam fsm_init = 0;
  wire [35-1:0] padr_0;
  wire [20-1:0] padr_bits_1;
  assign padr_bits_1 = 0;
  wire [29-1:0] truncR_2;
  wire [29-1:0] padl_3;
  wire [28-1:0] padl_bits_4;
  wire [1-1:0] toSInt_5;
  assign toSInt_5 = 0;
  wire [28-1:0] toSInt_imm_6;
  wire [27-1:0] const_7;
  assign const_7 = 27'd55364812;
  assign toSInt_imm_6 = { toSInt_5, const_7 };
  assign padl_bits_4 = toSInt_imm_6;
  assign padl_3 = { { 1{ padl_bits_4[27] } }, padl_bits_4 };
  assign truncR_2 = padl_3;
  wire [15-1:0] truncR_shift_8;
  assign truncR_shift_8 = truncR_2 >>> 14;
  wire [15-1:0] truncR_imm_9;
  assign truncR_imm_9 = (truncR_2[28])? truncR_shift_8[14:0] : truncR_2[28:14];
  assign padr_0 = { truncR_imm_9, padr_bits_1 };
  wire [13-1:0] truncR_10;
  wire [14-1:0] truncval_11;
  wire [15-1:0] toUsInt_12;
  wire [35-1:0] truncR_13;
  assign truncR_13 = o;
  wire [15-1:0] truncR_shift_14;
  assign truncR_shift_14 = truncR_13 >>> 20;
  wire [15-1:0] truncR_imm_15;
  assign truncR_imm_15 = (truncR_13[34])? truncR_shift_14[14:0] : truncR_13[34:20];
  assign toUsInt_12 = truncR_imm_15;
  assign truncval_11 = toUsInt_12[11:0];
  assign truncR_10 = truncval_11[12:0];
  wire [32-1:0] padl_16;
  wire [18-1:0] padl_bits_17;
  wire [33-1:0] truncR_18;
  wire [33-1:0] padl_19;
  wire [17-1:0] padl_bits_20;
  wire [95-1:0] truncR_21;
  wire [163-1:0] truncval_22;
  wire [163-1:0] padl_23;
  wire [85-1:0] padl_bits_24;
  wire [85-1:0] padl_25;
  wire [52-1:0] padl_bits_26;
  wire [98-1:0] truncR_27;
  wire [105-1:0] truncval_28;
  wire [105-1:0] padl_29;
  wire [52-1:0] padl_bits_30;
  wire [52-1:0] padr_31;
  wire [41-1:0] padr_bits_32;
  assign padr_bits_32 = 0;
  wire [1-1:0] toSInt_33;
  assign toSInt_33 = 0;
  wire [11-1:0] toSInt_imm_34;
  assign toSInt_imm_34 = { toSInt_33, n };
  assign padr_31 = { toSInt_imm_34, padr_bits_32 };
  assign padl_bits_30 = padr_31;
  assign padl_29 = { { 53{ padl_bits_30[51] } }, padl_bits_30 };
  wire [105-1:0] padl_35;
  wire [52-1:0] padl_bits_36;
  wire [52-1:0] padl_37;
  wire [50-1:0] padl_bits_38;
  wire [50-1:0] param_39;
  assign param_39 = n_to_response_time;
  assign padl_bits_38 = param_39;
  assign padl_37 = { { 2{ padl_bits_38[49] } }, padl_bits_38 };
  assign padl_bits_36 = padl_37;
  assign padl_35 = { { 53{ padl_bits_36[51] } }, padl_bits_36 };
  assign truncval_28 = padl_29 * padl_35;
  wire [98-1:0] truncval_imm_40;
  assign truncval_imm_40 = { truncval_28[104], truncval_28[96:0] };
  assign truncR_27 = truncval_imm_40;
  wire [52-1:0] truncR_shift_41;
  assign truncR_shift_41 = truncR_27 >>> 46;
  wire [52-1:0] truncR_imm_42;
  assign truncR_imm_42 = (truncR_27[97])? truncR_shift_41[51:0] : truncR_27[97:46];
  wire [52-1:0] padr_43;
  wire [2-1:0] padr_bits_44;
  assign padr_bits_44 = 0;
  wire [94-1:0] truncR_45;
  wire [101-1:0] truncval_46;
  wire [101-1:0] padl_47;
  wire [50-1:0] padl_bits_48;
  wire [50-1:0] padr_49;
  wire [39-1:0] padr_bits_50;
  assign padr_bits_50 = 0;
  wire [1-1:0] toSInt_51;
  assign toSInt_51 = 0;
  wire [11-1:0] toSInt_imm_52;
  assign toSInt_imm_52 = { toSInt_51, p };
  assign padr_49 = { toSInt_imm_52, padr_bits_50 };
  assign padl_bits_48 = padr_49;
  assign padl_47 = { { 51{ padl_bits_48[49] } }, padl_bits_48 };
  wire [101-1:0] padl_53;
  wire [50-1:0] padl_bits_54;
  wire [50-1:0] padl_55;
  wire [48-1:0] padl_bits_56;
  wire [48-1:0] param_57;
  assign param_57 = p_to_response_time;
  assign padl_bits_56 = param_57;
  assign padl_55 = { { 2{ padl_bits_56[47] } }, padl_bits_56 };
  assign padl_bits_54 = padl_55;
  assign padl_53 = { { 51{ padl_bits_54[49] } }, padl_bits_54 };
  assign truncval_46 = padl_47 * padl_53;
  wire [94-1:0] truncval_imm_58;
  assign truncval_imm_58 = { truncval_46[100], truncval_46[92:0] };
  assign truncR_45 = truncval_imm_58;
  wire [50-1:0] truncR_shift_59;
  assign truncR_shift_59 = truncR_45 >>> 44;
  wire [50-1:0] truncR_imm_60;
  assign truncR_imm_60 = (truncR_45[93])? truncR_shift_59[49:0] : truncR_45[93:44];
  assign padr_43 = { truncR_imm_60, padr_bits_44 };
  wire [52-1:0] padr_61;
  wire [8-1:0] padr_bits_62;
  assign padr_bits_62 = 0;
  wire [44-1:0] padl_63;
  wire [43-1:0] padl_bits_64;
  wire [1-1:0] toSInt_65;
  assign toSInt_65 = 0;
  wire [43-1:0] toSInt_imm_66;
  wire [42-1:0] param_67;
  assign param_67 = const_response_time;
  assign toSInt_imm_66 = { toSInt_65, param_67 };
  assign padl_bits_64 = toSInt_imm_66;
  assign padl_63 = { { 1{ padl_bits_64[42] } }, padl_bits_64 };
  assign padr_61 = { padl_63, padr_bits_62 };
  assign padl_bits_26 = truncR_imm_42 + padr_43 + padr_61;
  assign padl_25 = { { 33{ padl_bits_26[51] } }, padl_bits_26 };
  assign padl_bits_24 = padl_25;
  assign padl_23 = { { 78{ padl_bits_24[84] } }, padl_bits_24 };
  wire [163-1:0] padl_68;
  wire [85-1:0] padl_bits_69;
  wire [85-1:0] padr_70;
  wire [50-1:0] padr_bits_71;
  assign padr_bits_71 = 0;
  wire [1-1:0] toSInt_72;
  assign toSInt_72 = 0;
  wire [35-1:0] toSInt_imm_73;
  wire [34-1:0] const_74;
  assign const_74 = 34'd78125000;
  assign toSInt_imm_73 = { toSInt_72, const_74 };
  assign padr_70 = { toSInt_imm_73, padr_bits_71 };
  assign padl_bits_69 = padr_70;
  assign padl_68 = { { 78{ padl_bits_69[84] } }, padl_bits_69 };
  assign truncval_22 = padl_23 * padl_68;
  assign truncR_21 = truncval_22[94:0];
  assign padl_bits_20 = truncR_21[94:78];
  wire [16-1:0] padl_bits_zero_75;
  assign padl_bits_zero_75 = 0;
  assign padl_19 = { padl_bits_zero_75, padl_bits_20 };
  assign truncR_18 = padl_19;
  assign padl_bits_17 = truncR_18[32:15];
  wire [14-1:0] padl_bits_zero_76;
  assign padl_bits_zero_76 = 0;
  assign padl_16 = { padl_bits_zero_76, padl_bits_17 };
  assign wait_time = padl_16;
  wire [35-1:0] padr_77;
  wire [20-1:0] padr_bits_78;
  assign padr_bits_78 = 0;
  wire [29-1:0] truncR_79;
  wire [29-1:0] padl_80;
  wire [28-1:0] padl_bits_81;
  wire [1-1:0] toSInt_82;
  assign toSInt_82 = 0;
  wire [28-1:0] toSInt_imm_83;
  wire [27-1:0] const_84;
  assign const_84 = 27'd55364812;
  assign toSInt_imm_83 = { toSInt_82, const_84 };
  assign padl_bits_81 = toSInt_imm_83;
  assign padl_80 = { { 1{ padl_bits_81[27] } }, padl_bits_81 };
  assign truncR_79 = padl_80;
  wire [15-1:0] truncR_shift_85;
  assign truncR_shift_85 = truncR_79 >>> 14;
  wire [15-1:0] truncR_imm_86;
  assign truncR_imm_86 = (truncR_79[28])? truncR_shift_85[14:0] : truncR_79[28:14];
  assign padr_77 = { truncR_imm_86, padr_bits_78 };
  wire [13-1:0] truncR_87;
  wire [14-1:0] truncval_88;
  wire [15-1:0] toUsInt_89;
  wire [35-1:0] truncR_90;
  assign truncR_90 = o;
  wire [15-1:0] truncR_shift_91;
  assign truncR_shift_91 = truncR_90 >>> 20;
  wire [15-1:0] truncR_imm_92;
  assign truncR_imm_92 = (truncR_90[34])? truncR_shift_91[14:0] : truncR_90[34:20];
  assign toUsInt_89 = truncR_imm_92;
  assign truncval_88 = toUsInt_89[11:0];
  assign truncR_87 = truncval_88[12:0];
  wire [51-1:0] padr_93;
  wire [6-1:0] padr_bits_94;
  assign padr_bits_94 = 0;
  wire [46-1:0] truncval_95;
  wire [47-1:0] toUsInt_96;
  wire [88-1:0] truncR_97;
  wire [95-1:0] truncval_98;
  wire [95-1:0] padl_99;
  wire [47-1:0] padl_bits_100;
  wire [47-1:0] padr_101;
  wire [36-1:0] padr_bits_102;
  assign padr_bits_102 = 0;
  wire [1-1:0] toSInt_103;
  assign toSInt_103 = 0;
  wire [11-1:0] toSInt_imm_104;
  assign toSInt_imm_104 = { toSInt_103, n };
  assign padr_101 = { toSInt_imm_104, padr_bits_102 };
  assign padl_bits_100 = padr_101;
  assign padl_99 = { { 48{ padl_bits_100[46] } }, padl_bits_100 };
  wire [95-1:0] padl_105;
  wire [47-1:0] padl_bits_106;
  wire [47-1:0] padl_107;
  wire [45-1:0] padl_bits_108;
  wire [45-1:0] param_109;
  assign param_109 = n_to_tau;
  assign padl_bits_108 = param_109;
  assign padl_107 = { { 2{ padl_bits_108[44] } }, padl_bits_108 };
  assign padl_bits_106 = padl_107;
  assign padl_105 = { { 48{ padl_bits_106[46] } }, padl_bits_106 };
  assign truncval_98 = padl_99 * padl_105;
  wire [88-1:0] truncval_imm_110;
  assign truncval_imm_110 = { truncval_98[94], truncval_98[86:0] };
  assign truncR_97 = truncval_imm_110;
  wire [47-1:0] truncR_shift_111;
  assign truncR_shift_111 = truncR_97 >>> 41;
  wire [47-1:0] truncR_imm_112;
  assign truncR_imm_112 = (truncR_97[87])? truncR_shift_111[46:0] : truncR_97[87:41];
  wire [47-1:0] padl_113;
  wire [46-1:0] padl_bits_114;
  wire [1-1:0] toSInt_115;
  assign toSInt_115 = 0;
  wire [46-1:0] toSInt_imm_116;
  wire [86-1:0] truncR_117;
  wire [92-1:0] truncval_118;
  wire [92-1:0] padl_119;
  wire [46-1:0] padl_bits_120;
  wire [46-1:0] padr_121;
  wire [36-1:0] padr_bits_122;
  assign padr_bits_122 = 0;
  assign padr_121 = { p, padr_bits_122 };
  assign padl_bits_120 = padr_121;
  wire [46-1:0] padl_bits_zero_123;
  assign padl_bits_zero_123 = 0;
  assign padl_119 = { padl_bits_zero_123, padl_bits_120 };
  wire [92-1:0] padl_124;
  wire [46-1:0] padl_bits_125;
  wire [46-1:0] padl_126;
  wire [43-1:0] padl_bits_127;
  wire [43-1:0] param_128;
  assign param_128 = p_to_tau;
  assign padl_bits_127 = param_128;
  wire [3-1:0] padl_bits_zero_129;
  assign padl_bits_zero_129 = 0;
  assign padl_126 = { padl_bits_zero_129, padl_bits_127 };
  assign padl_bits_125 = padl_126;
  wire [46-1:0] padl_bits_zero_130;
  assign padl_bits_zero_130 = 0;
  assign padl_124 = { padl_bits_zero_130, padl_bits_125 };
  assign truncval_118 = padl_119 * padl_124;
  assign truncR_117 = truncval_118[85:0];
  assign toSInt_imm_116 = { toSInt_115, truncR_117[85:41] };
  assign padl_bits_114 = toSInt_imm_116;
  assign padl_113 = { { 1{ padl_bits_114[45] } }, padl_bits_114 };
  wire [47-1:0] padr_131;
  wire [4-1:0] padr_bits_132;
  assign padr_bits_132 = 0;
  wire [43-1:0] padl_133;
  wire [42-1:0] padl_bits_134;
  wire [1-1:0] toSInt_135;
  assign toSInt_135 = 0;
  wire [42-1:0] toSInt_imm_136;
  wire [41-1:0] param_137;
  assign param_137 = const_tau;
  assign toSInt_imm_136 = { toSInt_135, param_137 };
  assign padl_bits_134 = toSInt_imm_136;
  assign padl_133 = { { 1{ padl_bits_134[41] } }, padl_bits_134 };
  assign padr_131 = { padl_133, padr_bits_132 };
  assign toUsInt_96 = truncR_imm_112 + padl_113 + padr_131;
  assign truncval_95 = toUsInt_96[43:0];
  assign padr_93 = { truncval_95[44:0], padr_bits_94 };
  assign tau = padr_93;
  wire [13-1:0] truncR_138;
  wire [14-1:0] truncval_139;
  wire [15-1:0] toUsInt_140;
  wire [35-1:0] truncR_141;
  assign truncR_141 = o;
  wire [15-1:0] truncR_shift_142;
  assign truncR_shift_142 = truncR_141 >>> 20;
  wire [15-1:0] truncR_imm_143;
  assign truncR_imm_143 = (truncR_141[34])? truncR_shift_142[14:0] : truncR_141[34:20];
  assign toUsInt_140 = truncR_imm_143;
  assign truncval_139 = toUsInt_140[11:0];
  assign truncR_138 = truncval_139[12:0];
  wire [36-1:0] padl_144;
  wire [13-1:0] padl_bits_145;
  wire [36-1:0] truncR_146;
  wire [60-1:0] truncR_147;
  wire [93-1:0] truncval_148;
  wire [93-1:0] padl_149;
  wire [46-1:0] padl_bits_150;
  wire [46-1:0] padl_151;
  wire [16-1:0] padl_bits_152;
  wire [16-1:0] neg_imm_153;
  wire [16-1:0] padr_154;
  wire [2-1:0] padr_bits_155;
  assign padr_bits_155 = 0;
  wire [15-1:0] truncval_156;
  wire [35-1:0] truncR_157;
  assign truncR_157 = o;
  wire [15-1:0] truncR_shift_158;
  assign truncR_shift_158 = truncR_157 >>> 20;
  wire [15-1:0] truncR_imm_159;
  assign truncR_imm_159 = (truncR_157[34])? truncR_shift_158[14:0] : truncR_157[34:20];
  assign truncval_156 = truncR_imm_159;
  wire [14-1:0] truncval_imm_160;
  assign truncval_imm_160 = { truncval_156[14], truncval_156[12:0] };
  assign padr_154 = { truncval_imm_160, padr_bits_155 };
  assign neg_imm_153 = -padr_154;
  assign padl_bits_152 = neg_imm_153;
  assign padl_151 = { { 30{ padl_bits_152[15] } }, padl_bits_152 };
  assign padl_bits_150 = padl_151;
  assign padl_149 = { { 47{ padl_bits_150[45] } }, padl_bits_150 };
  wire [93-1:0] padl_161;
  wire [46-1:0] padl_bits_162;
  wire [46-1:0] padr_163;
  wire [12-1:0] padr_bits_164;
  assign padr_bits_164 = 0;
  wire [1-1:0] toSInt_165;
  assign toSInt_165 = 0;
  wire [34-1:0] toSInt_imm_166;
  wire [51-1:0] truncval_167;
  assign truncval_167 = 52'd2251799813685248 / tau;
  assign toSInt_imm_166 = { toSInt_165, truncval_167[32:0] };
  assign padr_163 = { toSInt_imm_166, padr_bits_164 };
  assign padl_bits_162 = padr_163;
  assign padl_161 = { { 47{ padl_bits_162[45] } }, padl_bits_162 };
  assign truncval_148 = padl_149 * padl_161;
  wire [60-1:0] truncval_imm_168;
  assign truncval_imm_168 = { truncval_148[92], truncval_148[58:0] };
  assign truncR_147 = truncval_imm_168;
  wire [36-1:0] truncR_shift_169;
  assign truncR_shift_169 = truncR_147 >>> 24;
  wire [36-1:0] truncR_imm_170;
  assign truncR_imm_170 = (truncR_147[59])? truncR_shift_169[35:0] : truncR_147[59:24];
  assign truncR_146 = truncR_imm_170;
  wire [13-1:0] truncR_shift_171;
  assign truncR_shift_171 = truncR_146 >>> 23;
  wire [13-1:0] truncR_imm_172;
  assign truncR_imm_172 = (truncR_146[35])? truncR_shift_171[12:0] : truncR_146[35:23];
  assign padl_bits_145 = truncR_imm_172;
  assign padl_144 = { { 23{ padl_bits_145[12] } }, padl_bits_145 };
  assign dvdt = padl_144;
  wire [35-1:0] padr_173;
  wire [20-1:0] padr_bits_174;
  assign padr_bits_174 = 0;
  wire [19-1:0] truncR_175;
  wire [19-1:0] padl_176;
  wire [16-1:0] padl_bits_177;
  wire [97-1:0] truncR_178;
  wire [168-1:0] truncval_179;
  wire [168-1:0] padl_180;
  wire [95-1:0] padl_bits_181;
  wire [95-1:0] padl_182;
  wire [60-1:0] padl_bits_183;
  wire [1-1:0] toSInt_184;
  assign toSInt_184 = 0;
  wire [60-1:0] toSInt_imm_185;
  wire [59-1:0] const_186;
  assign const_186 = 59'd57646075;
  assign toSInt_imm_185 = { toSInt_184, const_186 };
  assign padl_bits_183 = toSInt_imm_185;
  assign padl_182 = { { 35{ padl_bits_183[59] } }, padl_bits_183 };
  assign padl_bits_181 = padl_182;
  assign padl_180 = { { 73{ padl_bits_181[94] } }, padl_bits_181 };
  wire [168-1:0] padl_187;
  wire [95-1:0] padl_bits_188;
  wire [95-1:0] padr_189;
  wire [59-1:0] padr_bits_190;
  assign padr_bits_190 = 0;
  assign padr_189 = { dvdt, padr_bits_190 };
  assign padl_bits_188 = padr_189;
  assign padl_187 = { { 73{ padl_bits_188[94] } }, padl_bits_188 };
  assign truncval_179 = padl_180 * padl_187;
  wire [97-1:0] truncval_imm_191;
  assign truncval_imm_191 = { truncval_179[167], truncval_179[95:0] };
  assign truncR_178 = truncval_imm_191;
  wire [16-1:0] truncR_shift_192;
  assign truncR_shift_192 = truncR_178 >>> 81;
  wire [16-1:0] truncR_imm_193;
  assign truncR_imm_193 = (truncR_178[96])? truncR_shift_192[15:0] : truncR_178[96:81];
  assign padl_bits_177 = truncR_imm_193;
  assign padl_176 = { { 3{ padl_bits_177[15] } }, padl_bits_177 };
  assign truncR_175 = padl_176;
  wire [15-1:0] truncR_shift_194;
  assign truncR_shift_194 = truncR_175 >>> 4;
  wire [15-1:0] truncR_imm_195;
  assign truncR_imm_195 = (truncR_175[18])? truncR_shift_194[14:0] : truncR_175[18:4];
  assign padr_173 = { truncR_imm_195, padr_bits_174 };
  wire [32-1:0] padl_196;
  wire [2-1:0] padl_bits_197;
  wire [13-1:0] truncR_198;
  wire [17-1:0] truncR_199;
  wire [17-1:0] padl_200;
  wire [16-1:0] padl_bits_201;
  wire [92-1:0] truncR_202;
  wire [161-1:0] truncval_203;
  wire [161-1:0] padl_204;
  wire [84-1:0] padl_bits_205;
  wire [84-1:0] padl_206;
  wire [51-1:0] padl_bits_207;
  wire [98-1:0] truncR_208;
  wire [105-1:0] truncval_209;
  wire [105-1:0] padl_210;
  wire [52-1:0] padl_bits_211;
  wire [52-1:0] padr_212;
  wire [41-1:0] padr_bits_213;
  assign padr_bits_213 = 0;
  wire [1-1:0] toSInt_214;
  assign toSInt_214 = 0;
  wire [11-1:0] toSInt_imm_215;
  assign toSInt_imm_215 = { toSInt_214, n };
  assign padr_212 = { toSInt_imm_215, padr_bits_213 };
  assign padl_bits_211 = padr_212;
  assign padl_210 = { { 53{ padl_bits_211[51] } }, padl_bits_211 };
  wire [105-1:0] padl_216;
  wire [52-1:0] padl_bits_217;
  wire [52-1:0] padl_218;
  wire [50-1:0] padl_bits_219;
  wire [50-1:0] param_220;
  assign param_220 = n_to_response_time_lh;
  assign padl_bits_219 = param_220;
  assign padl_218 = { { 2{ padl_bits_219[49] } }, padl_bits_219 };
  assign padl_bits_217 = padl_218;
  assign padl_216 = { { 53{ padl_bits_217[51] } }, padl_bits_217 };
  assign truncval_209 = padl_210 * padl_216;
  wire [98-1:0] truncval_imm_221;
  assign truncval_imm_221 = { truncval_209[104], truncval_209[96:0] };
  assign truncR_208 = truncval_imm_221;
  wire [51-1:0] truncR_shift_222;
  assign truncR_shift_222 = truncR_208 >>> 47;
  wire [51-1:0] truncR_imm_223;
  assign truncR_imm_223 = (truncR_208[97])? truncR_shift_222[50:0] : truncR_208[97:47];
  wire [51-1:0] padr_224;
  wire [1-1:0] padr_bits_225;
  assign padr_bits_225 = 0;
  wire [94-1:0] truncR_226;
  wire [101-1:0] truncval_227;
  wire [101-1:0] padl_228;
  wire [50-1:0] padl_bits_229;
  wire [50-1:0] padr_230;
  wire [39-1:0] padr_bits_231;
  assign padr_bits_231 = 0;
  wire [1-1:0] toSInt_232;
  assign toSInt_232 = 0;
  wire [11-1:0] toSInt_imm_233;
  assign toSInt_imm_233 = { toSInt_232, p };
  assign padr_230 = { toSInt_imm_233, padr_bits_231 };
  assign padl_bits_229 = padr_230;
  assign padl_228 = { { 51{ padl_bits_229[49] } }, padl_bits_229 };
  wire [101-1:0] padl_234;
  wire [50-1:0] padl_bits_235;
  wire [50-1:0] padl_236;
  wire [48-1:0] padl_bits_237;
  wire [48-1:0] param_238;
  assign param_238 = p_to_response_time_lh;
  assign padl_bits_237 = param_238;
  assign padl_236 = { { 2{ padl_bits_237[47] } }, padl_bits_237 };
  assign padl_bits_235 = padl_236;
  assign padl_234 = { { 51{ padl_bits_235[49] } }, padl_bits_235 };
  assign truncval_227 = padl_228 * padl_234;
  wire [94-1:0] truncval_imm_239;
  assign truncval_imm_239 = { truncval_227[100], truncval_227[92:0] };
  assign truncR_226 = truncval_imm_239;
  wire [50-1:0] truncR_shift_240;
  assign truncR_shift_240 = truncR_226 >>> 44;
  wire [50-1:0] truncR_imm_241;
  assign truncR_imm_241 = (truncR_226[93])? truncR_shift_240[49:0] : truncR_226[93:44];
  assign padr_224 = { truncR_imm_241, padr_bits_225 };
  wire [51-1:0] padr_242;
  wire [6-1:0] padr_bits_243;
  assign padr_bits_243 = 0;
  wire [45-1:0] padl_244;
  wire [44-1:0] padl_bits_245;
  wire [1-1:0] toSInt_246;
  assign toSInt_246 = 0;
  wire [44-1:0] toSInt_imm_247;
  wire [43-1:0] param_248;
  assign param_248 = const_response_time_lh;
  assign toSInt_imm_247 = { toSInt_246, param_248 };
  assign padl_bits_245 = toSInt_imm_247;
  assign padl_244 = { { 1{ padl_bits_245[43] } }, padl_bits_245 };
  assign padr_242 = { padl_244, padr_bits_243 };
  assign padl_bits_207 = truncR_imm_223 + padr_224 + padr_242;
  assign padl_206 = { { 33{ padl_bits_207[50] } }, padl_bits_207 };
  assign padl_bits_205 = padl_206;
  assign padl_204 = { { 77{ padl_bits_205[83] } }, padl_bits_205 };
  wire [161-1:0] padl_249;
  wire [84-1:0] padl_bits_250;
  wire [84-1:0] padr_251;
  wire [49-1:0] padr_bits_252;
  assign padr_bits_252 = 0;
  wire [1-1:0] toSInt_253;
  assign toSInt_253 = 0;
  wire [35-1:0] toSInt_imm_254;
  wire [34-1:0] const_255;
  assign const_255 = 34'd78125000;
  assign toSInt_imm_254 = { toSInt_253, const_255 };
  assign padr_251 = { toSInt_imm_254, padr_bits_252 };
  assign padl_bits_250 = padr_251;
  assign padl_249 = { { 77{ padl_bits_250[83] } }, padl_bits_250 };
  assign truncval_203 = padl_204 * padl_249;
  assign truncR_202 = truncval_203[91:0];
  assign padl_bits_201 = truncR_202[91:76];
  wire [1-1:0] padl_bits_zero_256;
  assign padl_bits_zero_256 = 0;
  assign padl_200 = { padl_bits_zero_256, padl_bits_201 };
  assign truncR_199 = padl_200;
  assign truncR_198 = truncR_199[16:4];
  assign padl_bits_197 = truncR_198[12:11];
  wire [30-1:0] padl_bits_zero_257;
  assign padl_bits_zero_257 = 0;
  assign padl_196 = { padl_bits_zero_257, padl_bits_197 };
  assign wait_time_lh = padl_196;
  wire [35-1:0] padr_258;
  wire [20-1:0] padr_bits_259;
  assign padr_bits_259 = 0;
  wire [41-1:0] truncR_260;
  wire [41-1:0] padl_261;
  wire [37-1:0] padl_bits_262;
  wire [1-1:0] toSInt_263;
  assign toSInt_263 = 0;
  wire [37-1:0] toSInt_imm_264;
  wire [36-1:0] const_265;
  assign const_265 = 36'd68719476;
  assign toSInt_imm_264 = { toSInt_263, const_265 };
  assign padl_bits_262 = toSInt_imm_264;
  assign padl_261 = { { 4{ padl_bits_262[36] } }, padl_bits_262 };
  assign truncR_260 = padl_261;
  wire [15-1:0] truncR_shift_266;
  assign truncR_shift_266 = truncR_260 >>> 26;
  wire [15-1:0] truncR_imm_267;
  assign truncR_imm_267 = (truncR_260[40])? truncR_shift_266[14:0] : truncR_260[40:26];
  assign padr_258 = { truncR_imm_267, padr_bits_259 };
  wire [13-1:0] truncR_268;
  wire [14-1:0] truncval_269;
  wire [15-1:0] toUsInt_270;
  wire [35-1:0] truncR_271;
  assign truncR_271 = o;
  wire [15-1:0] truncR_shift_272;
  assign truncR_shift_272 = truncR_271 >>> 20;
  wire [15-1:0] truncR_imm_273;
  assign truncR_imm_273 = (truncR_271[34])? truncR_shift_272[14:0] : truncR_271[34:20];
  assign toUsInt_270 = truncR_imm_273;
  assign truncval_269 = toUsInt_270[11:0];
  assign truncR_268 = truncval_269[12:0];
  wire [59-1:0] padr_274;
  wire [10-1:0] padr_bits_275;
  assign padr_bits_275 = 0;
  wire [50-1:0] truncval_276;
  wire [51-1:0] toUsInt_277;
  wire [51-1:0] padr_278;
  wire [3-1:0] padr_bits_279;
  assign padr_bits_279 = 0;
  wire [48-1:0] padl_280;
  wire [47-1:0] padl_bits_281;
  wire [1-1:0] toSInt_282;
  assign toSInt_282 = 0;
  wire [47-1:0] toSInt_imm_283;
  wire [88-1:0] truncR_284;
  wire [94-1:0] truncval_285;
  wire [94-1:0] padl_286;
  wire [47-1:0] padl_bits_287;
  wire [47-1:0] padr_288;
  wire [37-1:0] padr_bits_289;
  assign padr_bits_289 = 0;
  assign padr_288 = { n, padr_bits_289 };
  assign padl_bits_287 = padr_288;
  wire [47-1:0] padl_bits_zero_290;
  assign padl_bits_zero_290 = 0;
  assign padl_286 = { padl_bits_zero_290, padl_bits_287 };
  wire [94-1:0] padl_291;
  wire [47-1:0] padl_bits_292;
  wire [47-1:0] padl_293;
  wire [44-1:0] padl_bits_294;
  wire [44-1:0] param_295;
  assign param_295 = n_to_tau_lh;
  assign padl_bits_294 = param_295;
  wire [3-1:0] padl_bits_zero_296;
  assign padl_bits_zero_296 = 0;
  assign padl_293 = { padl_bits_zero_296, padl_bits_294 };
  assign padl_bits_292 = padl_293;
  wire [47-1:0] padl_bits_zero_297;
  assign padl_bits_zero_297 = 0;
  assign padl_291 = { padl_bits_zero_297, padl_bits_292 };
  assign truncval_285 = padl_286 * padl_291;
  assign truncR_284 = truncval_285[87:0];
  assign toSInt_imm_283 = { toSInt_282, truncR_284[87:42] };
  assign padl_bits_281 = toSInt_imm_283;
  assign padl_280 = { { 1{ padl_bits_281[46] } }, padl_bits_281 };
  assign padr_278 = { padl_280, padr_bits_279 };
  wire [96-1:0] truncR_298;
  wire [103-1:0] truncval_299;
  wire [103-1:0] padl_300;
  wire [51-1:0] padl_bits_301;
  wire [51-1:0] padr_302;
  wire [40-1:0] padr_bits_303;
  assign padr_bits_303 = 0;
  wire [1-1:0] toSInt_304;
  assign toSInt_304 = 0;
  wire [11-1:0] toSInt_imm_305;
  assign toSInt_imm_305 = { toSInt_304, p };
  assign padr_302 = { toSInt_imm_305, padr_bits_303 };
  assign padl_bits_301 = padr_302;
  assign padl_300 = { { 52{ padl_bits_301[50] } }, padl_bits_301 };
  wire [103-1:0] padl_306;
  wire [51-1:0] padl_bits_307;
  wire [51-1:0] padl_308;
  wire [49-1:0] padl_bits_309;
  wire [49-1:0] param_310;
  assign param_310 = p_to_tau_lh;
  assign padl_bits_309 = param_310;
  assign padl_308 = { { 2{ padl_bits_309[48] } }, padl_bits_309 };
  assign padl_bits_307 = padl_308;
  assign padl_306 = { { 52{ padl_bits_307[50] } }, padl_bits_307 };
  assign truncval_299 = padl_300 * padl_306;
  wire [96-1:0] truncval_imm_311;
  assign truncval_imm_311 = { truncval_299[102], truncval_299[94:0] };
  assign truncR_298 = truncval_imm_311;
  wire [51-1:0] truncR_shift_312;
  assign truncR_shift_312 = truncR_298 >>> 45;
  wire [51-1:0] truncR_imm_313;
  assign truncR_imm_313 = (truncR_298[95])? truncR_shift_312[50:0] : truncR_298[95:45];
  wire [51-1:0] padr_314;
  wire [6-1:0] padr_bits_315;
  assign padr_bits_315 = 0;
  wire [45-1:0] padl_316;
  wire [44-1:0] padl_bits_317;
  wire [1-1:0] toSInt_318;
  assign toSInt_318 = 0;
  wire [44-1:0] toSInt_imm_319;
  wire [43-1:0] param_320;
  assign param_320 = const_tau_lh;
  assign toSInt_imm_319 = { toSInt_318, param_320 };
  assign padl_bits_317 = toSInt_imm_319;
  assign padl_316 = { { 1{ padl_bits_317[43] } }, padl_bits_317 };
  assign padr_314 = { padl_316, padr_bits_315 };
  assign toUsInt_277 = padr_278 + truncR_imm_313 + padr_314;
  assign truncval_276 = toUsInt_277[47:0];
  assign padr_274 = { truncval_276[48:0], padr_bits_275 };
  assign tau_lh = padr_274;
  wire [33-1:0] truncR_321;
  wire [34-1:0] truncval_322;
  wire [35-1:0] toUsInt_323;
  assign toUsInt_323 = o;
  assign truncval_322 = toUsInt_323[31:0];
  assign truncR_321 = truncval_322[32:0];
  wire [37-1:0] padl_324;
  wire [13-1:0] padl_bits_325;
  wire [37-1:0] truncR_326;
  wire [97-1:0] truncR_327;
  wire [131-1:0] truncval_328;
  wire [131-1:0] padl_329;
  wire [65-1:0] padl_bits_330;
  wire [65-1:0] padl_331;
  wire [35-1:0] padl_bits_332;
  wire [35-1:0] padr_333;
  wire [6-1:0] padr_bits_334;
  assign padr_bits_334 = 0;
  wire [29-1:0] padl_335;
  wire [28-1:0] padl_bits_336;
  wire [1-1:0] toSInt_337;
  assign toSInt_337 = 0;
  wire [28-1:0] toSInt_imm_338;
  wire [27-1:0] const_339;
  assign const_339 = 27'd55364812;
  assign toSInt_imm_338 = { toSInt_337, const_339 };
  assign padl_bits_336 = toSInt_imm_338;
  assign padl_335 = { { 1{ padl_bits_336[27] } }, padl_bits_336 };
  assign padr_333 = { padl_335, padr_bits_334 };
  assign padl_bits_332 = padr_333 - o;
  assign padl_331 = { { 30{ padl_bits_332[34] } }, padl_bits_332 };
  assign padl_bits_330 = padl_331;
  assign padl_329 = { { 66{ padl_bits_330[64] } }, padl_bits_330 };
  wire [131-1:0] padl_340;
  wire [65-1:0] padl_bits_341;
  wire [65-1:0] padr_342;
  wire [30-1:0] padr_bits_343;
  assign padr_bits_343 = 0;
  wire [1-1:0] toSInt_344;
  assign toSInt_344 = 0;
  wire [35-1:0] toSInt_imm_345;
  wire [59-1:0] truncval_346;
  assign truncval_346 = 60'd576460752303423488 / tau_lh;
  assign toSInt_imm_345 = { toSInt_344, truncval_346[33:0] };
  assign padr_342 = { toSInt_imm_345, padr_bits_343 };
  assign padl_bits_341 = padr_342;
  assign padl_340 = { { 66{ padl_bits_341[64] } }, padl_bits_341 };
  assign truncval_328 = padl_329 * padl_340;
  wire [97-1:0] truncval_imm_347;
  assign truncval_imm_347 = { truncval_328[130], truncval_328[95:0] };
  assign truncR_327 = truncval_imm_347;
  wire [37-1:0] truncR_shift_348;
  assign truncR_shift_348 = truncR_327 >>> 60;
  wire [37-1:0] truncR_imm_349;
  assign truncR_imm_349 = (truncR_327[96])? truncR_shift_348[36:0] : truncR_327[96:60];
  assign truncR_326 = truncR_imm_349;
  wire [13-1:0] truncR_shift_350;
  assign truncR_shift_350 = truncR_326 >>> 24;
  wire [13-1:0] truncR_imm_351;
  assign truncR_imm_351 = (truncR_326[36])? truncR_shift_350[12:0] : truncR_326[36:24];
  assign padl_bits_325 = truncR_imm_351;
  assign padl_324 = { { 24{ padl_bits_325[12] } }, padl_bits_325 };
  assign dodt = padl_324;
  wire [35-1:0] padr_352;
  wire [17-1:0] padr_bits_353;
  assign padr_bits_353 = 0;
  wire [18-1:0] padl_354;
  wire [17-1:0] padl_bits_355;
  wire [98-1:0] truncR_356;
  wire [169-1:0] truncval_357;
  wire [169-1:0] padl_358;
  wire [96-1:0] padl_bits_359;
  wire [96-1:0] padl_360;
  wire [60-1:0] padl_bits_361;
  wire [1-1:0] toSInt_362;
  assign toSInt_362 = 0;
  wire [60-1:0] toSInt_imm_363;
  wire [59-1:0] const_364;
  assign const_364 = 59'd57646075;
  assign toSInt_imm_363 = { toSInt_362, const_364 };
  assign padl_bits_361 = toSInt_imm_363;
  assign padl_360 = { { 36{ padl_bits_361[59] } }, padl_bits_361 };
  assign padl_bits_359 = padl_360;
  assign padl_358 = { { 73{ padl_bits_359[95] } }, padl_bits_359 };
  wire [169-1:0] padl_365;
  wire [96-1:0] padl_bits_366;
  wire [96-1:0] padr_367;
  wire [59-1:0] padr_bits_368;
  assign padr_bits_368 = 0;
  assign padr_367 = { dodt, padr_bits_368 };
  assign padl_bits_366 = padr_367;
  assign padl_365 = { { 73{ padl_bits_366[95] } }, padl_bits_366 };
  assign truncval_357 = padl_358 * padl_365;
  wire [98-1:0] truncval_imm_369;
  assign truncval_imm_369 = { truncval_357[168], truncval_357[96:0] };
  assign truncR_356 = truncval_imm_369;
  wire [17-1:0] truncR_shift_370;
  assign truncR_shift_370 = truncR_356 >>> 81;
  wire [17-1:0] truncR_imm_371;
  assign truncR_imm_371 = (truncR_356[97])? truncR_shift_370[16:0] : truncR_356[97:81];
  assign padl_bits_355 = truncR_imm_371;
  assign padl_354 = { { 1{ padl_bits_355[16] } }, padl_bits_355 };
  assign padr_352 = { padl_354, padr_bits_353 };
  assign out = (fsm == 0)? truncR_10[12:3] : truncR_87[12:3];

  always @(posedge clk) begin
    prev_sys_clk <= sys_clk;
  end

  localparam fsm_1 = 1;
  localparam fsm_2 = 2;
  localparam fsm_3 = 3;
  localparam fsm_4 = 4;

  always @(posedge clk) begin
    if(reset) begin
      fsm <= fsm_init;
    end else begin
      case(fsm)
        fsm_init: begin
          if(reset) begin
            o <= 35'd3543348019;
          end else begin
            o <= padr_0;
          end
          if(~prev_sys_clk & sys_clk & ((n > p) & (n <= 10'd512))) begin
            fsm <= fsm_1;
          end 
        end
        fsm_1: begin
          if(reset) begin
            o <= 35'd3543348019;
          end else begin
            o <= padr_77;
          end
          if(state_cycle_counter > wait_time) begin
            state_cycle_counter <= 0;
          end else begin
            state_cycle_counter <= state_cycle_counter + 1;
          end
          if(state_cycle_counter > wait_time) begin
            fsm <= fsm_2;
          end 
        end
        fsm_2: begin
          if(reset) begin
            o <= 35'd3543348019;
          end else begin
            o <= o + padr_173;
          end
          if(prev_sys_clk & ~sys_clk) begin
            fsm <= fsm_3;
          end 
        end
        fsm_3: begin
          if(reset) begin
            o <= 35'd3543348019;
          end else begin
            o <= padr_258;
          end
          if(state_cycle_counter > wait_time_lh) begin
            state_cycle_counter <= 0;
          end else begin
            state_cycle_counter <= state_cycle_counter + 1;
          end
          if(state_cycle_counter > wait_time_lh) begin
            fsm <= fsm_4;
          end 
        end
        fsm_4: begin
          if(reset) begin
            o <= 35'd3543348019;
          end else begin
            o <= o + padr_352;
          end
          if((o > 35'd3532610600) & (o <= 35'd17179869184)) begin
            fsm <= fsm_init;
          end 
        end
      endcase
    end
  end


endmodule

