`include "./sar_adc.v"
module stub;

sar_adc sar_inst();
endmodule